
library ieee;
use ieee.std_logic_1164.all;

entity logic_unit is
    port(
        a  : in  std_logic_vector(31 downto 0);
        b  : in  std_logic_vector(31 downto 0);
        op : in  std_logic_vector(1 downto 0);
        r  : out std_logic_vector(31 downto 0)
    );
end logic_unit;

architecture synth of logic_unit is
	signal result : std_logic_vector(31 downto 0);
begin
	checkOP : process (op, a, b)
	begin
		case op is
		when "00" => result <= a nor b;
		when "01" => result <= a and b;
		when "10" => result <= a or b;
		when "11" => result <= a xor b;
		when others => result <= (others => '0');
		end case; 
	end process CheckOP;
r <= result;
end synth;
